module main